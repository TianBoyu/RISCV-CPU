//the wb module have been down at the regfile.v